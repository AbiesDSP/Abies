module ${module_name} (
    input wire clk
);

endmodule
