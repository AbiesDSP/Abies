`timescale 1ns/1ps

module ${module_name} (
    input wire clk
);

endmodule
