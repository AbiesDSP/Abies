module ${module_name} (
    input logic clk
);

endmodule
