`default_nettype none

module ${module_name} (
    input wire clk
);

endmodule
